module top (in1,out);
input   in1;
output  out;

buf(out, in1);
endmodule
